*** Inversor ***

*parametros
.param SUPPLY=1.5
*.option scale=25n
.options savecurrents

*.nodeset V(1)=1.5

.temp 70

* fuentes
Vdd 1 0 'SUPPLY'
Vin 3 0 PULSE 0 'SUPPLY' (50ps 0ps 0ps 100ps 200ps)

* inversor
Mn1 4 3 0 0 tipoN
Mp1 4 3 1 1 tipoP


* Carga
*Cload 4 0 50n
Cload 0 4 50n

.model tipoN NMOS (LEVEL=3 PHI=0.600000 TOX=2.1500E-08 XJ=0.200000U TPG=1 VTO=0.8063 DELTA=9.4090E-01 LD=1.3540E-07 KP=1.0877E-04 UO=680.4 THETA=8.3620E-02 RSH=109.3 GAMMA=0.5487 NSUB=2.3180E+16 NFS=1.98E+12 VMAX=1.8700E+05 ETA=5.5740E-02 KAPPA=5.9210E-02 CGDO=3.2469E-10 CGSO=3.2469E-10 CGBO=3.7124E-10 CJ=3.1786E-04 MJ=1.0148 CJSW=1.3284E-10 MJSW=0.119521 PB=0.800000)
.model tipoP PMOS (LEVEL=3 PHI=0.600000 TOX=2.1500E-08 XJ=0.200000U TPG=-1 VTO=-0.9403 DELTA=8.5790E-01LD=1.1650E-09 KP=3.4276E-05 UO=214.4 THETA=1.4010E-01 RSH=122.2 GAMMA=0.5615 NSUB=2.4270E+16 NFS=3.46E+12 VMAX=3.9310E+05 ETA=1.5670E-01 KAPPA=9.9990E+00 CGDO=2.7937E-12 CGSO=2.7937E-12 CGBO=3.5981E-10 CJ=4.5952E-04 MJ=0.4845 CJSW=2.7917E-10 MJSW=0.365250 PB=0.850000)

*.model tipoN NMOS (W=4 L=2 AS=20 PS=18 AD=20 PD=18)
*.model tipoP PMOS (W=8 L=2 AS=40 PS=26 AD=40 PD=26)


.tran 1ps 1ns UIC

.control
run

*plotting
plot v(4)
plot v(3)
plot v(3) v(4)
plot @Cload[i]
*plot @Cload[i] vs v(3)

.endc

.end
