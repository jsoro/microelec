*
* Test of MOS BSIM3 implementation; DC transfer curve
****************************************************************** 
MN1 13 2 0 4 NMOS 
MN2 23 2 0 5 NMOS 
MN3 33 2 0 6 NMOS   
MN4 43 2 0 7 NMOS   
MN5 53 2 0 8 NMOS 
** L=10U W=50.0U AD=100P AS=100P PD=40U PS=40U 
VDS 3 0 0.05    
VGS 2 0 0
V1 3 13 0       
V2 3 23 0       
V3 3 33 0       
V4 3 43 0       
V5 3 53 0       
VBS1 4 0 0      
VBS2 5 0 -1
VBS3 6 0 -2     
VBS4 7 0 -3
VBS5 8 0 -4     
*************************************************************** 
.OPTIONS LIMPTS=5000 ACCT       
.DC VGS 0 5 0.01
.PRINT DC I(V1) I(V2) I(V3) I(V4) I(V5) 
*.PLOT DC I(V1) I(V2) I(V3) I(V4) I(V5) 
*.OPTIONS LIMPTS=501 ACCT       
*VGS  2  0  PWL(0 0 5 5)
*.TRAN 0 5 0.01
*.PRINT TRAN I(V1) I(V2) I(V3) I(V4) I(V5) 
***** MODEL PARAMETERS TEMP3 ********************       
* This file contains the BSIM3 process file parameters as they should
* be input to the .model card of spice3c1.
.model NMOS  nmos level=8
+ Tnom=27.0
+ nch= 1.024685E+17  tox=1.00000E-08 xj=1.00000E-07
+ lint= 3.75860E-08 wint=-2.02101528644562E-07
+ vth0= .6094574   k1= .5341038  k2= 1.703463E-03  k3=-17.24589
+ dvt0= .1767506  dvt1= .5109418  dvt2=-0.05
+ nlx= 9.979638E-08  w0=1e-6
+ k3b= 4.139039
+ vsat= 97662.05  ua=-1.748481E-09  ub= 3.178541E-18  uc=1.3623e-10 
+ rdsw= 298.873  u0= 307.2991 prwb=-2.24e-4
+ a0= .4976366
+ keta=-2.195445E-02  a1= .0332883  a2= .9
+ voff=-9.623903E-02  nFactor= .8408191  cit= 3.994609E-04
+ cdsc= 1.130797E-04
+ cdscb=2.4e-5
+ eta0= .0145072  etab=-3.870303E-03
+ dsub= .4116711
+ pclm= 1.813153  pdiblc1= 2.003703E-02  pdiblc2= .00129051 pdiblcb=-1.034e-3
+ drout= .4380235  pscbe1= 5.752058E+08  pscbe2= 7.510319E-05
+ pvag= .6370527 prt=68.7 ngate=1.e20 alpha0=1.e-7 beta0=28.4 
+ prwg=-0.001 ags=1.2
+ dvt0w=0.58 dvt1w=5.3e6 dvt2w=-0.0032
+ kt1=-.3  kt2=-.03
+ at= 33000
+ ute=-1.5
+ ua1= 4.31E-09  ub1= 7.61E-18  uc1=-2.378e-10
+ kt1l=1e-8
+ wr=1 b0=1e-7 b1=1e-7 dwg=5e-8 dwb=2e-8 delta=0.015
+ cgdl=1e-10 cgsl=1e-10 cgbo=1e-10 xpart=0.0
+ cgdo=0.4e-9 cgso=0.4e-9 
+ clc=0.1e-6
+ cle=0.6
+ ckappa=0.6


.model PMOS  pmos level=8
+ Tnom=27.0
+ nch= 5.73068E+16  tox=1.00000E-08 xj=1.00000E-07
+ lint= 8.195860E-08 wint=-1.821562E-07
+ vth0= -.86094574   k1= .341038  k2= 2.703463E-02  k3=12.24589
+ dvt0= .767506  dvt1= .65109418  dvt2=-0.145
+ nlx= 1.979638E-07  w0=1.1e-6
+ k3b= -2.4139039
+ vsat= 60362.05  ua=1.348481E-09  ub= 3.178541E-19  uc=1.1623e-10 
+ rdsw= 498.873  u0= 137.2991 prwb=-1.2e-5
+ a0= .3276366
+ keta=-1.8195445E-02  a1= .0232883  a2= .9
+ voff=-6.623903E-02  nFactor= 1.0408191  cit= 4.994609E-04
+ cdsc= 1.030797E-3
+ cdscb=2.84e-4
+ eta0= .0245072  etab=-1.570303E-03
+ dsub= .24116711
+ pclm= 2.6813153  pdiblc1= 4.003703E-02  pdiblc2= .00329051 pdiblcb=-2.e-4
+ drout= .1380235  pscbe1= 0  pscbe2=1.e-28 
+ pvag= -.16370527
+ prwg=-0.001 ags=1.2
+ dvt0w=0.58 dvt1w=5.3e6 dvt2w=-0.0032
+ kt1=-.3  kt2=-.03 prt=76.4
+ at= 33000
+ ute=-1.5
+ ua1= 4.31E-09  ub1= 7.61E-18  uc1=-2.378e-10
+ kt1l=0
+ wr=1 b0=1e-7 b1=1e-7 dwg=5e-8 dwb=2e-8 delta=0.015
+ cgdl=1e-10 cgsl=1e-10 cgbo=1e-10 xpart=0.0
+ cgdo=0.4e-9 cgso=0.4e-9 
+ clc=0.1e-6
+ cle=0.6
+ ckappa=0.6
.END
