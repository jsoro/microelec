*** Inversor ***

*parametros
.param SUPPLY=4.20
*.option scale=25n
.options savecurrents



.temp 70

* fuentes
Vdd 1 0 'SUPPLY'
Vin 3 0 PULSE 0 'SUPPLY' (50ps 0ps 0ps 100ps 200ps)

* inversor
Mn1 4 3 0 0 tipoN
Mp1 4 3 1 1 tipoP


* Carga

*Cload 4 0 50n
Cload 0 4 50n

.model tipoN NMOS (LEVEL=3 PHI=0.600000 TOX=2.1200E-08 XJ=0.200000U TPG=1 VTO=0.7860 DELTA=6.9670E-01 LD=1.6470E-07 KP=9.6379E-05 UO=591.7 THETA=8.1220E-02 RSH=8.5450E+01 GAMMA=0.5863 NSUB=2.7470E+16 NFS=1.98E+12 VMAX=1.7330E+05 ETA=4.3680E-02 KAPPA=1.3960E-01 CGDO=4.0241E-10 CGSO=4.0241E-10 CGBO=3.6144E-10 CJ=3.8541E MJ=0.5027 CJSW=1.6457E-10 MJSW=0.217168 PB=0.850000)

.model tipoP PMOS (LEVEL=3 PHI=0.600000 TOX=2.1200E-08 XJ=0.200000U TPG=-1 VTO=-0.9056 DELTA=1.5200E+00 LD=2.2000E-08 KP=2.9352E-05 UO=180.2 THETA=1.2480E-01 RSH=1.0470E+02 GAMMA=0.4863 NSUB=1.8900E+16 NFS=3.46E+12 VMAX=3.7320E+05 ETA=1.6410E-01 KAPPA=9.6940E+00 CGDO=5.3752E-11 CGSO=5.3752E-11 CGBO=3.3650E-10 CJ=4.8447E-04 MJ=0.5027 CJSW=1.6457E-10 MJSW=0.217168 PB=0.850000)

*.model tipoN NMOS (W=4 L=2 AS=20 PS=18 AD=20 PD=18)
*.model tipoP PMOS (W=8 L=2 AS=40 PS=26 AD=40 PD=26)


.tran 1ps 1ns

.control
run

*plotting
plot v(4)
plot v(3)
plot v(3) v(4)
plot @Cload[i]
*plot @Cload[i] vs v(3)

*.endc

.end
