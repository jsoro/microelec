NetListTina (TINA Netlist Editor format)
**************************************
**  This file was created by TINA   **
**         www.tina.com             ** 
**      (c) DesignSoft, Inc.        **          
**     www.designsoftware.com       **
**************************************
.LIB "<TINADIR>\EXAMPLES\SPICE\TSPICE.LIB"
.LIB "<TINADIR>\SPICELIB\Operational Amplifiers.LIB"
.TEMP 27
.AC DEC 20 10 1MEG
.TRAN 400U 200M UIC
.DC LIN VG3 0 1 10M

.PROBE V(3,0)

VG3         1 4 DC 0 AC 1 0
+ PWL TIME_SCALE_FACTOR=20M VALUE_SCALE_FACTOR=5
+      REPEAT FOREVER
+       (0, 0) (50N 1) (499.99995M 1) (500.00005M -1) (999.99995M -1) (1,0) ENDREPEAT
VG3_DC      4 0 5
VG4         2 0 DC 0 AC 1 0
+ PULSE ( 0 5 0  0  0  1e19 1e20 )
MT3         2 1 3 3  ME_2N6804_P_1 NRD=0 NRS=0 
MT4         3 1 0 0  ME_2N6755_N_1 NRD=0 NRS=0 
C2          3 0 1U 

.MODEL ME_2N6804_P_1 PMOS( LEVEL=3 VTO=-3.695 KP=10.41U PHI=600M GAMMA=0 TOX=100N 
+      UO=300 VMAX=0 DELTA=0 THETA=0 ETA=0 
+      L=2U W=1.2 RD=66.52M RS=153M RG=4.931 
+      RB=0 RDS=444.4MEG IS=5.483P N=3 PB=800M 
+      CBD=1.291N CBS=0 MJ=500M TT=295N CGSO=1.783N 
+      CGDO=134.9P CGBO=0 KF=0 AF=1 )
.MODEL ME_2N6755_N_1 NMOS( LEVEL=3 VTO=3.128 KP=21.14U PHI=600M GAMMA=0 TOX=100N 
+      UO=600 VMAX=0 DELTA=0 THETA=0 ETA=0 
+      L=2U W=1.1 RD=64.68M RS=120.7M RG=5.839 
+      RB=0 RDS=600K IS=44.14F N=1 PB=800M 
+      CBD=1.261N CBS=0 MJ=500M TT=370N CGSO=725.6P 
+      CGDO=310.6P CGBO=0 KF=0 AF=1 )

.END
