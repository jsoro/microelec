*** SPICE deck for cell NOR3{lay} from library inversor
*** Created on Wed Jun 03, 2020 17:04:27
*** Last revised on Tue Jun 09, 2020 16:42:30
*** Written on Tue Jun 09, 2020 16:44:06 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NOR3{lay}
Mnmos@0 Y B gnd gnd N L=0.4U W=1U AS=5.84P AD=3.18P PS=15.2U PD=10.8U
Mnmos@1 Y C gnd gnd N L=0.4U W=1U AS=5.84P AD=3.18P PS=15.2U PD=10.8U
Mnmos@2 Y A gnd gnd N L=0.4U W=1U AS=5.84P AD=3.18P PS=15.2U PD=10.8U
Mpmos@0 net@3 B net@2 vdd P L=0.4U W=2U AS=5.56P AD=5.78P PS=11.2U PD=9.6U
Mpmos@1 Y C net@3 vdd P L=0.4U W=2U AS=5.78P AD=3.18P PS=9.6U PD=10.8U
Mpmos@2 net@2 A vdd vdd P L=0.4U W=2U AS=15.56P AD=5.56P PS=37.2U PD=11.2U

* Spice Code nodes in cell cell 'NOR3{lay}'
vdd VDD 0 DC 5
vinA A 0 pulse 0 5 0 1n 1n .5m 1m
vinB B 0 pulse 0 5 0 1n 1n .2m 1m
vinC C 0 pulse 0 5 0 1n 3n .2m .5m
.tran 0 2m
.END
