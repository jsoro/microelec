*** SPICE deck for cell AOI22{lay} from library tarea5
*** Created on Wed Jun 03, 2020 17:04:27
*** Last revised on Tue Jun 09, 2020 18:19:26
*** Written on Sat Jun 13, 2020 11:24:04 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: AOI22{lay}
Mnmos@0 gnd B net@0 gnd N L=0.4U W=1U AS=3.16P AD=10.14P PS=8.6U PD=24.8U
Mnmos@1 net@24 C Y gnd N L=0.4U W=1U AS=2.67P AD=3.01P PS=8.7U PD=7.9U
Mnmos@2 net@0 A Y gnd N L=0.4U W=1U AS=2.67P AD=3.16P PS=8.7U PD=8.6U
Mnmos@3 gnd D net@24 gnd N L=0.4U W=1U AS=3.01P AD=10.14P PS=7.9U PD=24.8U
Mpmos@0 Y B net@2 vdd P L=0.4U W=2U AS=3.74P AD=2.67P PS=11.8U PD=8.7U
Mpmos@1 net@2 C vdd vdd P L=0.4U W=2U AS=19.2P AD=3.74P PS=25.2U PD=11.8U
Mpmos@2 Y A net@2 vdd P L=0.4U W=2U AS=3.74P AD=2.67P PS=11.8U PD=8.7U
Mpmos@3 net@2 D vdd vdd P L=0.4U W=2U AS=19.2P AD=3.74P PS=25.2U PD=11.8U

* Spice Code nodes in cell cell 'AOI22{lay}'
vdd VDD 0 DC 5
vinA A 0 pulse 0 5 0 1n 1n .5m 1m
vinB B 0 pulse 0 5 0 1n 1n .2m 1m
vinC C 0 pulse 0 5 0 1n 3n .2m .5m
vinD D 0 pulse 0 5 0 1n 3n .1m .3m
.tran 0 2m
.END
