*** SPICE deck for cell NAND3{lay} from library inversor
*** Created on Wed Jun 03, 2020 17:04:27
*** Last revised on Tue Jun 09, 2020 16:21:07
*** Written on Tue Jun 09, 2020 16:28:21 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND3{lay}
Mnmos@0 net@1 B net@0 gnd N L=0.4U W=1U AS=3.16P AD=2.88P PS=8.6U PD=7.4U
Mnmos@1 Y C net@1 gnd N L=0.4U W=1U AS=2.88P AD=3.34P PS=7.4U PD=10.8U
Mnmos@2 net@0 A gnd gnd N L=0.4U W=1U AS=13.96P AD=3.16P PS=33.2U PD=8.6U
Mpmos@0 Y B vdd vdd P L=0.4U W=2U AS=7.44P AD=3.34P PS=18.533U PD=10.8U
Mpmos@1 Y C vdd vdd P L=0.4U W=2U AS=7.44P AD=3.34P PS=18.533U PD=10.8U
Mpmos@2 Y A vdd vdd P L=0.4U W=2U AS=7.44P AD=3.34P PS=18.533U PD=10.8U

* Spice Code nodes in cell cell 'NAND3{lay}'
vdd VDD 0 DC 5
vinA A 0 pulse 0 5 0 1n 1n .5m 1m
vinB B 0 pulse 0 5 0 1n 1n .2m 1m
vinC C 0 pulse 0 5 0 1n 3n .2m .5m
.tran 0 2m
.END
