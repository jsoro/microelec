*** Inversor ***

*parametros
.param SUPPLY=1.5
*.option scale=25n
.options savecurrents

*.nodeset V(1)=1.5

.temp 70

* fuentes
Vdd 1 0 'SUPPLY'
Vin 3 0 PULSE 0 'SUPPLY' (50ps 0ps 0ps 100ps 200ps)

* inversor
Mn1 4 3 0 0 tipoN
Mp1 4 3 1 1 tipoP


* Carga
*Cload 4 0 50n
Cload 0 4 50n

.model tipoN NMOS (LEVEL=3 PHI=0.600000 TOX=2.0500E-08 XJ=0.200000U TPG=1 VTO=0.8147 DELTA=3.0170E-05 LD=1.7540E-07 KP=8.9765E-05 UO=532.9 THETA=9.0470E-02 RSH=1.5870E+01 GAMMA=0.6654 NSUB=3.7840E+16 NFS=5.5000E+12 VMAX=1.7140E+05 ETA=6.4550E-02 KAPPA=5.6190E-02 CGDO=4.4318E-10 CGSO=4.4318E-10 CGBO=3.2044E-10 CJ=3.1786E-04 MJ=1.0148 CJSW=1.3284E-10 MJSW=0.119521 PB=0.800000)
.model tipoP PMOS (LEVEL=3 PHI=0.600000 TOX=2.0500E-08 XJ=0.200000U TPG=-1 VTO=-0.9189 DELTA=2.3190E+00 LD=1.0440E-08 KP=3.3521E-05  UO=199.0 THETA=1.7940E-01 RSH=25.0000 GAMMA=0.4124 NSUB=1.4540E+16 NFS=5.0000E+12 VMAX=5.4640E+05 ETA=2.1090E-01 KAPPA=9.3670E+00 CGDO=2.6379E-11 CGSO=2.6379E-11 CGBO=2.8996E-10 CJ=4.6135E-04 MJ=0.4831 CJSW=1.8681E-10 MJSW=0.315030 PB=0.850000)

*.model tipoN NMOS (W=4 L=2 AS=20 PS=18 AD=20 PD=18)
*.model tipoP PMOS (W=8 L=2 AS=40 PS=26 AD=40 PD=26)


.tran 1ps 1ns UIC

.control
run

*plotting
plot v(4)
plot v(3)
plot v(3) v(4)
plot @Cload[i]
*plot @Cload[i] vs v(3)

.endc

.end
