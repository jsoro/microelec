* First line is ignored

*** SUBCIRCUIT layout_inversor FROM CELL layout_inversor{lay}
.SUBCKT layout_inversor 0 A vdd Y
Mnmos_0 Y A 0 0 N L=0.4U W=1U
Mpmos_0 Y A vdd vdd P L=0.4U W=2U
.ENDS layout_inversor
